CIRCUIT C:\microwind2\Book on CMOS\ChargePump.MSK
*
* IC Technology: CMOS 0.12�m - 6 Metal
*
VDD 1 0 DC 1.20
Vclock1 8 0 PULSE(0.00 1.20 0.50N 0.05N 0.05N 0.50N 1.10N)
*
* List of nodes
* "VCharge" corresponds to n�4
* "N5" corresponds to n�5
* "Vout" corresponds to n�6
* "clock1" corresponds to n�8
* "N9" corresponds to n�9
*
* MOS devices
MN1 4 4 6 0 N1  W= 0.60U L= 0.12U
MN2 0 8 5 0 N1  W= 0.36U L= 0.12U
MP1 4 4 1 1 P1  W= 0.60U L= 0.12U
MP2 1 8 5 1 P1  W= 0.96U L= 0.12U
*
C2 1 0  2.540fF
C3 1 0  1.250fF
C4 4 0 17.788fF
C5 5 0 17.199fF
C6 6 0  0.705fF
C8 8 0  0.660fF
C9 9 0  0.119fF
*
* Crosstalk capacitance
*
Cx4_5 4 5 1.305fF
Cx5_9 5 9 0.108fF
*
* n-MOS Model 3 :
* low leakage
.MODEL N1 NMOS LEVEL=3 VTO=0.40 U0=0.060 TOX= 3.0E-9
+LD =0.000U THETA=0.300 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=170.00K
+CGSO=  0.0p CGDO=  0.0p
* high speed
.MODEL N2 NMOS LEVEL=3 VTO=0.30 U0=0.060 TOX= 3.0E-9
+LD =0.000U THETA=0.300 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=170.00K
+CGSO=  0.0p CGDO=  0.0p
* high voltage
.MODEL N3 NMOS LEVEL=3 VTO=0.70 U0=0.060 TOX= 7.0E-9
+LD =0.000U THETA=0.300 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=170.00K
+CGSO=  0.0p CGDO=  0.0p
*
* p-MOS Model 3:
* high speed pMOS
.MODEL P1 PMOS LEVEL=3 VTO=-0.40 U0=0.020 TOX= 3.0E-9
+LD =0.000U THETA=0.300 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=120.00K
+CGSO=  0.0p CGDO=  0.0p
* high speed
.MODEL P2 PMOS LEVEL=3 VTO=-0.30 U0=0.020 TOX= 3.0E-9
+LD =0.000U THETA=0.300 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=120.00K
+CGSO=  0.0p CGDO=  0.0p
* high voltage
.MODEL P3 PMOS LEVEL=3 VTO=-0.70 U0=0.020 TOX= 7.0E-9
+LD =0.000U THETA=0.300 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=120.00K
+CGSO=  0.0p CGDO=  0.0p
*
* Transient analysis
*
.TEMP 27.0
.TRAN 0.30PS 10.00N
.PROBE
.END
